
module SB_RAM256x16
  #(parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000)
   (
    output [15:0] RDATA,
    input         RCLK,
    input         RCLKE,
    input         RE,
    input [7:0]   RADDR,
    input         WCLK,
    input         WCLKE,
    input         WE,
    input [7:0]   WADDR,
    input [15:0]  MASK,
    input [15:0]  WDATA
    );

   SB_RAM40_4K #(.INIT_0(INIT_0),
                 .INIT_1(INIT_1),
                 .INIT_2(INIT_2),
                 .INIT_3(INIT_3),
                 .INIT_4(INIT_4),
                 .INIT_5(INIT_5),
                 .INIT_6(INIT_6),
                 .INIT_7(INIT_7),
                 .INIT_8(INIT_8),
                 .INIT_9(INIT_9),
                 .INIT_A(INIT_A),
                 .INIT_B(INIT_B),
                 .INIT_C(INIT_C),
                 .INIT_D(INIT_D),
                 .INIT_E(INIT_E),
                 .INIT_F(INIT_F))
   u_ram40_4k (.RDATA(RDATA),
               .RADDR(RADDR),
               .RCLK(RCLK),
               .RCLKE(RCLKE),
               .RE(RE),
               .WADDR(WADDR),
               .WCLK(WCLK),
               .WCLKE(WCLKE),
               .WDATA(WDATA),
               .WE(WE),
               .MASK(MASK));
endmodule
